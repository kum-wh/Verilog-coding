`timescale 1ns / 1ps
//actually does the loading screen
module frame(input clock, [12:0] index, output reg ennd = 0 , reg [15:0] data );
    reg [24:0] COUNT = 25'b0;
    reg [2:0] COUNT2 = 3'b0;
    always @ (posedge clock) begin
        COUNT <= COUNT + 1;
        COUNT2 <= (COUNT == 25'b0)?COUNT2 + 1:COUNT2;
        ennd <= (COUNT2 == 3'b111)?1:ennd;
       
        case(COUNT2)
        3'b000: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=24)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=24)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=24)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=24)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b001: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=32)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=32)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=32)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=32)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b010: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=40)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=40)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=40)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=40)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b011: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=48)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=48)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=48)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=48)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b100: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=56)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=56)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=56)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=56)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b101: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=64)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=64)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=64)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=64)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b110: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=72)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=72)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=72)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=72)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        3'b111: data <= (index/96==24)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==38)?16'b1111111111111111:(index%96==39)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==48)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==60)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==25)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==54)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==26)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==27)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:16'b0):
                        (index/96==28)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==43)?16'b1111111111111111:(index%96==44)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==55)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==61)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==29)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==30)?((index%96==33)?16'b1111111111111111:(index%96==37)?16'b1111111111111111:(index%96==40)?16'b1111111111111111:(index%96==42)?16'b1111111111111111:(index%96==45)?16'b1111111111111111:(index%96==47)?16'b1111111111111111:(index%96==49)?16'b1111111111111111:(index%96==51)?16'b1111111111111111:(index%96==53)?16'b1111111111111111:(index%96==56)?16'b1111111111111111:(index%96==57)?16'b1111111111111111:(index%96==59)?16'b1111111111111111:(index%96==62)?16'b1111111111111111:16'b0):
                        (index/96==31)?((index%96<32)?16'b0:(index%96>62)?16'b0:(index%96==36)?16'b0:(index%96==41)?16'b0:(index%96==43)?16'b0:(index%96==44)?16'b0:(index%96==46)?16'b0:(index%96==49)?16'b0:(index%96==50)?16'b0:(index%96==52)?16'b0:(index%96==54)?16'b0:(index%96==55)?16'b0:(index%96==58)?16'b0:16'b1111111111111111):
                        (index/96==35)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):
                        (index/96==36)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=78)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==37)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=78)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==38)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=78)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==39)?((index%96==16)?16'b1111111111111111:(index%96==79)?16'b1111111111111111:((index%96>=17)?((index%96<=78)?16'b0000000000011111:16'b0):16'b0)):
                        (index/96==40)?((index%96<16)?16'b0:(index%96>79)?16'b0:16'b1111111111111111):16'b0;
        endcase
    end
endmodule
